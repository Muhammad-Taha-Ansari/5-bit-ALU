module multiplier(input [4:0] A, input [4:0] B, output [9:0] product);
    assign product = A * B;
endmodule
