module Shift_Left(input [4:0] A, output [4:0] shifted);
    assign shifted = A << 1;
endmodule
